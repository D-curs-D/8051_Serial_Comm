.title KiCad schematic
IC1 EN RW RS NC_01 NC_02 MOSI MISO SCK RESET Rx Tx Net-_IC1-Pad12_ NC_03 NC_04 NC_05 NC_06 NC_07 XTAL2 XTAL1 GND DATA7 DATA6 DATA5 DATA4 DATA3 DATA2 DATA1 DATA0 NC_08 NC_09 Vin NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 Vin AT89S52-24PU
C3 Vin RESET 10uF
R1 RESET GND 10k
U1 VCC GND Vin1 LM7805_TO220
C1 VCC GND 100nF
C5 Vin1 GND 10nF
D4 Vin1 GND 1N4007
D2 Vin Vin1 1N5818
D3 Vin Vin2 1N5818
SW1 RESET Vin SW_SPST
SW2 GND Net-_IC1-Pad12_ SW_SPST
Y1 XTAL2 XTAL1 Crystal_Small
P1 MOSI Vin2 SCK MISO RESET GND CONN_02X03
D6 GND Rx LED_Small
D7 GND Tx LED_Small
R2 VCC Net-_D1-Pad2_ 330
D1 GND Net-_D1-Pad2_ Blue
J1 Net-_D5-Pad1_ GND Screw_Terminal_01x02
D5 Net-_D5-Pad1_ VCC 1N4007
J2 Rx Tx Conn_02x01
R3 Net-_DS1-Pad16_ GND 220
RV1 NC_18 Net-_DS1-Pad3_ GND 10k
C2 XTAL2 GND 22pF
C4 XTAL1 GND 22pF
J3 GND Vin1 Net-_DS1-Pad3_ RS RW EN DATA0 DATA1 DATA2 DATA3 DATA4 DATA5 DATA6 DATA7 Vin1 Net-_DS1-Pad16_ Conn_01x16_Female
DS1 GND Vin1 Net-_DS1-Pad3_ RS RW EN DATA0 DATA1 DATA2 DATA3 DATA4 DATA5 DATA6 DATA7 Vin1 Net-_DS1-Pad16_ WC1602A
.end
